package test_pkg;
import uvm_pkg::*;
	`include "uvm_macros.svh"
	//`include "tb_defs.sv"
	`include "master_xtns.sv"
	`include "master_config.sv"
	`include "slave_config.sv"
	`include "env_config.sv"
	`include "master_seqs.sv"
	`include "master_seqr.sv"
	`include "master_mon.sv"
	`include "master_driver.sv"

	`include "master_agent.sv"
	`include "master_atop.sv"
	`include "slave_xtns.sv"
	`include "slave_mon.sv"
	`include "slave_seqr.sv"
	`include "slave_driver.sv"
	`include "slave_agent.sv"
	`include "slave_atop.sv"
	`include "score_board.sv"

	`include "tb.sv"


	`include "vtest.sv"
endpackage


